// partition.cdl
netcdf partition {
dimensions:
        P = 1 ;
        L = 1 ;
        NX = 30 ;
        NY = 30 ;

group: bounding_boxes {
  variables:
        int domain_x(P) ;
        int domain_y(P) ;
        int domain_extent_x(P) ;
        int domain_extent_y(P) ;
  data:

   domain_x = 0 ;

   domain_y = 0 ;

   domain_extent_x = 30 ;

   domain_extent_y = 30 ;
  } // group bounding_boxes
}

