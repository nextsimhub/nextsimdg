netcdf partition_metadata_2 {
dimensions:
	NX = 10 ;
	NY = 9 ;
	P = 2 ;
	T = 1 ;
	B = 1 ;
	L = UNLIMITED ; // (0 currently)
	R = UNLIMITED ; // (0 currently)

group: bounding_boxes {
  variables:
  	int domain_x(P) ;
  	int domain_y(P) ;
  	int domain_extent_x(P) ;
  	int domain_extent_y(P) ;
  data:

   domain_x = 0, 4 ;

   domain_y = 0, 0 ;

   domain_extent_x = 4, 6 ;

   domain_extent_y = 9, 9 ;
  } // group bounding_boxes

group: connectivity {
  variables:
  	int top_neighbors(P) ;
  	int top_neighbor_ids(T) ;
  	int top_neighbor_halos(T) ;
  	int bottom_neighbors(P) ;
  	int bottom_neighbor_ids(B) ;
  	int bottom_neighbor_halos(B) ;
  	int left_neighbors(P) ;
  	int left_neighbor_ids(L) ;
  	int left_neighbor_halos(L) ;
  	int right_neighbors(P) ;
  	int right_neighbor_ids(R) ;
  	int right_neighbor_halos(R) ;
  data:

   top_neighbors = 0, 1 ;

   top_neighbor_ids = 0 ;

   top_neighbor_halos = 9 ;

   bottom_neighbors = 1, 0 ;

   bottom_neighbor_ids = 1 ;

   bottom_neighbor_halos = 9 ;

   left_neighbors = 0, 0 ;

   right_neighbors = 0, 0 ;
  } // group connectivity
}
